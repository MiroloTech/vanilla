module project

pub struct Project {
	pub mut:
	path                  string
	hidden_file_pahts     []string
	name                  string
	run_command           string
}
