module ui

pub enum TextAlign {
	start
	centre
	end
}
