module ui

pub struct RenderInfo {
	pub mut:
	delta            f64
}
